`define ADDR_TIM_RCV_CORE_PHASE_MEAS_CTL1 5'h0
`define TIM_RCV_CORE_PHASE_MEAS_CTL1_NAVG_OFFSET 0
`define TIM_RCV_CORE_PHASE_MEAS_CTL1_NAVG 32'hffffffff
`define ADDR_TIM_RCV_CORE_DMTD_A_CTL   5'h4
`define TIM_RCV_CORE_DMTD_A_CTL_DEGLITCHER_THRES_OFFSET 0
`define TIM_RCV_CORE_DMTD_A_CTL_DEGLITCHER_THRES 32'h0000ffff
`define TIM_RCV_CORE_DMTD_A_CTL_RESERVED1_OFFSET 16
`define TIM_RCV_CORE_DMTD_A_CTL_RESERVED1 32'hffff0000
`define ADDR_TIM_RCV_CORE_DMTD_B_CTL   5'h8
`define TIM_RCV_CORE_DMTD_B_CTL_DEGLITCHER_THRES_OFFSET 0
`define TIM_RCV_CORE_DMTD_B_CTL_DEGLITCHER_THRES 32'h0000ffff
`define TIM_RCV_CORE_DMTD_B_CTL_RESERVED1_OFFSET 16
`define TIM_RCV_CORE_DMTD_B_CTL_RESERVED1 32'hffff0000
`define ADDR_TIM_RCV_CORE_PHASE_MEAS   5'hc
`define TIM_RCV_CORE_PHASE_MEAS_VAL_OFFSET 0
`define TIM_RCV_CORE_PHASE_MEAS_VAL 32'hffffffff
`define ADDR_TIM_RCV_CORE_F_DMTD_A     5'h10
`define TIM_RCV_CORE_F_DMTD_A_FREQ_OFFSET 0
`define TIM_RCV_CORE_F_DMTD_A_FREQ 32'h0fffffff
`define TIM_RCV_CORE_F_DMTD_A_VALID_OFFSET 28
`define TIM_RCV_CORE_F_DMTD_A_VALID 32'h10000000
`define ADDR_TIM_RCV_CORE_F_DMTD_B     5'h14
`define TIM_RCV_CORE_F_DMTD_B_FREQ_OFFSET 0
`define TIM_RCV_CORE_F_DMTD_B_FREQ 32'h0fffffff
`define TIM_RCV_CORE_F_DMTD_B_VALID_OFFSET 28
`define TIM_RCV_CORE_F_DMTD_B_VALID 32'h10000000
