`define ADDR_TIM_RCV_CORE_PHASE_MEAS_CTL1 4'h0
`define TIM_RCV_CORE_PHASE_MEAS_CTL1_NAVG_OFFSET 0
`define TIM_RCV_CORE_PHASE_MEAS_CTL1_NAVG 32'hffffffff
`define ADDR_TIM_RCV_CORE_DMTD_A_CTL   4'h4
`define TIM_RCV_CORE_DMTD_A_CTL_DEGLITCHER_THRES_OFFSET 0
`define TIM_RCV_CORE_DMTD_A_CTL_DEGLITCHER_THRES 32'h0000ffff
`define TIM_RCV_CORE_DMTD_A_CTL_RESERVED1_OFFSET 16
`define TIM_RCV_CORE_DMTD_A_CTL_RESERVED1 32'hffff0000
`define ADDR_TIM_RCV_CORE_DMTD_B_CTL   4'h8
`define TIM_RCV_CORE_DMTD_B_CTL_DEGLITCHER_THRES_OFFSET 0
`define TIM_RCV_CORE_DMTD_B_CTL_DEGLITCHER_THRES 32'h0000ffff
`define TIM_RCV_CORE_DMTD_B_CTL_RESERVED1_OFFSET 16
`define TIM_RCV_CORE_DMTD_B_CTL_RESERVED1 32'hffff0000
